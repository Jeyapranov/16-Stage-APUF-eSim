* C:\FOSSEE_2.3\eSim\library\SubcircuitLibrary\buffer\buffer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 1/29/2026 11:51:54 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad1_ /in Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M1  Net-_M1-Pad1_ /in GND GND mosfet_n		
M4  /out Net-_M1-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M3  /out Net-_M1-Pad1_ GND GND mosfet_n		
v2  Net-_M2-Pad3_ GND DC		
U1  /in /out PORT		

.end
